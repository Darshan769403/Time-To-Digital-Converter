**Time to Digital Converter**
.subckt inverter 1 2
m1 2 1 5 5 pmod l=1u w=100u
m2 2 1 0 0 nmod l=1u w=100
.model pmod pmos level=54 version=4.7
.model nmod nmos level=54 version=4.7
.ends
.subckt nand_gate 1 2 4
m1 3 2 0 0 nmod l=1u w=100u
m2 4 1 3 3 nmod l=1u w=100u
m3 4 1 5 5 pmod l=1u w=100u
m4 4 2 5 5 pmod l=1u w=100u
.model pmod pmos level=54 version=4.7
.model nmod nmos level=54 version=4.7
.ends
.subckt and_gate 1 2 6
m1 3 2 0 0 nmod l=1u w=100u
m2 4 1 3 3 nmod l=1u w=100u
m3 6 4 0 0 nmod l=1u w=100u
m4 4 1 5 5 pmod l=1u w=100u
m5 4 2 5 5 pmod l=1u w=100u
m6 6 4 5 5 pmod l=1u w=100u
.model pmod pmos level=54 version=4.7
.model nmod nmos level=54 version=4.7
.ends
.subckt dff 8 9 13 14
xa 8 10 inverter
xb 8 9 11 nand_gate
xc 9 10 12 nand_gate
xd 11 14 13 nand_gate
xe 13 12 14 nand_gate
.ends
Vdd 5 0 dc 5V
Vd1 20 0 pulse(0 5V 0 0 0 10ns 20ns)
Vd2 21 0 pulse(0 5V 0 0 0 10ns 50ns)
Vclk 22 0 pulse(0 5V 0 0 0 10ns 20ns)
xd1 20 22 23 24 dff
xd2 21 22 25 26 dff
xd1andd2 23 26 27 and_gate
xcounter 27 22 28 27 dff
.tran 0.1ns 60ns
.control
run
plot v(20) v(21)  v(28)
.endc
.end